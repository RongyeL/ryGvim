// +FHDR----------------------------------------------------------------------------
//                 Copyright (c) 2022 
//                       ALL RIGHTS RESERVED
// ---------------------------------------------------------------------------------
// Filename      : test.v
// Author        : Rongye
// Created On    : 2022-12-22 05:09
// Last Modified : 2022-12-22 05:13
// ---------------------------------------------------------------------------------
// Description   : 
//
//
// -FHDR----------------------------------------------------------------------------
module test (
    input   [3:0] clk,
    input           rst_n,
    output [4:0] data_o
    

);
    
endmodule

